// Section 3 
// Packages and the outermost structure of a bsv design

package TestPackage
    // TODO
endpackage