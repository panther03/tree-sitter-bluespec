x = 4 + 5;