ResultArbiter ra = test;